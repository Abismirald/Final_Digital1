library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity rom is
	port(
		cod_bcd: in std_logic_vector(3 downto 0); --es la salida del mux
		hc: in std_logic_vector(2 downto 0); -- bits 567
		vc: in std_logic_vector(2 downto 0); -- bits 567
		led: out std_logic		
		);
end;

architecture rom_arq of rom is

constant rom: std_logic_vector(0 to 767):= --767= 64(cada caracter)*12(cant caracteres) codificacion
"00111100"&"01111110"&"01100110"&"01100110"&"01100110"&"01100110"&"01111110"&"00111100"& --0 (0000)
"00011000"&"01111000"&"01111000"&"00011000"&"00011000"&"00011000"&"00011000"&"00011000"& --1 (0001)
"00111100"&"01111110"&"01100110"&"00001100"&"00011000"&"00110000"&"01111110"&"01111110"& --2 (0010)
"01111110"&"01111110"&"00001100"&"00011000"&"00001100"&"00000110"&"01111110"&"01111100"& --3 (0011)
"01100110"&"01100110"&"01100110"&"01111110"&"01111110"&"00000110"&"00000110"&"00000110"& --4 (0100)
"01111110"&"01111110"&"01100000"&"01111100"&"01111110"&"00000110"&"01111110"&"01111100"& --5 (0101)
"00001110"&"00011110"&"00110000"&"01100000"&"01111100"&"01100110"&"01111110"&"00111100"& --6 (0110)
"01111100"&"01111100"&"00001100"&"00111110"&"00111110"&"00001100"&"00001100"&"00001100"& --7 (0111)
"00111100"&"01111110"&"01100110"&"00111100"&"01111110"&"01100110"&"01111110"&"00111100"& --8 (1000)
"00111100"&"01111110"&"01100110"&"01111110"&"00111110"&"00000110"&"01111110"&"01111100"& --9 (1001)
"00000000"&"00000000"&"00000000"&"00000000"&"00000000"&"00000000"&"00011000"&"00011000"& --Punto(1010)
"01100110"&"01100110"&"01100110"&"01100110"&"01100110"&"00111100"&"00011000"&"00011000"; --V(1011)

signal cuenta: std_logic_vector(9 downto 0);
		
begin
	cuenta <= cod_bcd & vc & hc; 
	--la posicion estará dada por los 4b del bcd, los bit 567 del vc y los bit 567 del hc
	led <= rom(to_integer(unsigned(cuenta)));
end;